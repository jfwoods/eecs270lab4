module Calculator(KEY, SW, HEX7, HEX6, HEX5, HEX4, HEX3, HEX2, HEX0);
   input [2:0] KEY;
   input [7:0] SW; 
   output [6:0] HEX7, HEX6;
   output [6:0] HEX5, HEX4;
   output [6:0] HEX3, HEX2;
   output [6:0] HEX0; 

endmodule